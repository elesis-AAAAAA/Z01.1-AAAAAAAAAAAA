-- Elementos de Sistemas
-- by Luciano Soares
-- Ram8.vhd

Library ieee;
use ieee.std_logic_1164.all;

entity TopLevel is
	port(
		SW      : in  std_logic_vector(9 downto 0);
		LEDR     : out std_logic_vector(9 downto 0);
		KEY		 : in  std_logic_vector(3 downto 0);
		HEX0		: out std_logic_vector(6 downto 0);
		HEX1 : out std_logic_vector(6 downto 0);
		HEX2 : out std_logic_vector(6 downto 0);
		HEX3 : out std_logic_vector(6 downto 0)
	);
end entity;



architecture arch of TopLevel is

signal output_pc : std_logic_vector(15 downto 0);
signal input_pc : std_logic_vector(15 downto 0) := "0000000000000000";

component PC is
	port(
			clock     : in  STD_LOGIC;
			increment : in  STD_LOGIC;
			load      : in  STD_LOGIC;
			reset     : in  STD_LOGIC;
			input     : in  STD_LOGIC_VECTOR(15 downto 0);
			output    : out STD_LOGIC_VECTOR(15 downto 0)
	);
end component;

component sevenSeg is
	port (
			bcd : in  STD_LOGIC_VECTOR(3 downto 0);
			leds: out STD_LOGIC_VECTOR(6 downto 0));
end component;

begin


	pcpm: PC port map(
		clock => not KEY(0),
		increment => SW(0),
		load => SW(1),
		reset => SW(2),
		input => input_pc,
		output => output_pc
	);

	hex0port: sevenSeg port map (
		bcd => output_pc(3 downto 0),
		leds => HEX0);

	hex1port: sevenSeg port map (
		bcd => output_pc(7 downto 4),
		leds => HEX1);
	
	hex2port: sevenSeg port map (
		bcd => output_pc(11 downto 8),
		leds => HEX2);
	
	hex3port: sevenSeg port map (
		bcd => output_pc(15 downto 12),
		leds => HEX3);




end architecture;
